`include "cpu_data.v"

module CheckBranch(operator, check_branch, flags);

endmodule
